`include "CS_if.sv"

package CS_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "CS_transaction"
`include "CS_random_sequence.sv"
`include "CS_directed_sequence.sv"
`include "CS_sequencer.sv"
`include "CS_driver.sv"
`include "CS_monitor.sv"
`include "CS_scoreboard.sv"
`include "CS_agent.sv"
`include "CS_environment.sv"
`include "CS_base_test.sv"  
endpackage


